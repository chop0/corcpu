`timescale 1ns / 1ps

module frontend(

    );
endmodule

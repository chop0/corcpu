package instructions;
`define R_TYPE_INSTRUCTION(NAME, OPCODE, FUNCT3, FUNCT7) \
function [31:0] NAME(input [4:0] rd, rs1, rs2); \
    begin \
        NAME = {FUNCT7, rs2, rs1, FUNCT3, rd, OPCODE}; \
    end \
endfunction

// R-Type Instructions
`R_TYPE_INSTRUCTION(add, 7'b0110011, 3'b000, 7'b0000000)
`R_TYPE_INSTRUCTION(sub, 7'b0110011, 3'b000, 7'b0100000)
`R_TYPE_INSTRUCTION(xor_, 7'b0110011, 3'b100, 7'b0000000)
`R_TYPE_INSTRUCTION(or_, 7'b0110011, 3'b110, 7'b0000000)
`R_TYPE_INSTRUCTION(and_, 7'b0110011, 3'b111, 7'b0000000)
`R_TYPE_INSTRUCTION(sll, 7'b0110011, 3'b001, 7'b0000000)
`R_TYPE_INSTRUCTION(srl, 7'b0110011, 3'b101, 7'b0000000)
`R_TYPE_INSTRUCTION(sra, 7'b0110011, 3'b101, 7'b0100000)
`R_TYPE_INSTRUCTION(slt, 7'b0110011, 3'b010, 7'b0000000)
`R_TYPE_INSTRUCTION(sltu, 7'b0110011, 3'b011, 7'b0000000)

`define I_TYPE_INSTRUCTION(NAME, OPCODE, FUNCT3) \
function [31:0] NAME(input [4:0] rd, rs1, input [11:0] imm); \
    begin \
        NAME = {imm, rs1, FUNCT3, rd, OPCODE}; \
    end \
endfunction

// I-Type Instructions
`I_TYPE_INSTRUCTION(addi, 7'b0010011, 3'b000)
`I_TYPE_INSTRUCTION(xori, 7'b0010011, 3'b100)
`I_TYPE_INSTRUCTION(ori, 7'b0010011, 3'b110)
`I_TYPE_INSTRUCTION(andi, 7'b0010011, 3'b111)
`I_TYPE_INSTRUCTION(slli, 7'b0010011, 3'b001)
`I_TYPE_INSTRUCTION(srli, 7'b0010011, 3'b101)
`I_TYPE_INSTRUCTION(srai, 7'b0010011, 3'b101)
`I_TYPE_INSTRUCTION(slti, 7'b0010011, 3'b010)
`I_TYPE_INSTRUCTION(sltiu, 7'b0010011, 3'b011)

endpackage;
`ifndef CLASSES_SV
`define CLASSES_SV

package synchronous_fifo_tb;

endpackage

`endif